
module proj_qsys (
	clk_clk);	

	input		clk_clk;
endmodule
